-- Vhdl test bench created from schematic /home/luca/ISE_ws/FF_ms/ffms.sch - Thu Feb 21 19:36:27 2019
--
-- Notes: 
-- 1) This testbench template has been automatically generated using types
-- std_logic and std_logic_vector for the ports of the unit under test.
-- Xilinx recommends that these types always be used for the top-level
-- I/O of a design in order to guarantee that the testbench will bind
-- correctly to the timing (post-route) simulation model.
-- 2) To use this template as your testbench, change the filename to any
-- name of your choice with the extension .vhd, and use the "Source->Add"
-- menu in Project Navigator to import the testbench. Then
-- edit the user defined section below, adding code to generate the 
-- stimulus for your design.
--
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.numeric_std.ALL;
LIBRARY UNISIM;
USE UNISIM.Vcomponents.ALL;
ENTITY ffms_ffms_sch_tb IS
END ffms_ffms_sch_tb;
ARCHITECTURE behavioral OF ffms_ffms_sch_tb IS 

   COMPONENT ffms
   PORT( Clk	:	IN	STD_LOGIC; 
          D	:	IN	STD_LOGIC; 
          Q	:	OUT	STD_LOGIC);
   END COMPONENT;

   SIGNAL Clk	:	STD_LOGIC;
   SIGNAL D	:	STD_LOGIC;
   SIGNAL Q	:	STD_LOGIC;


constant Clk_period : time := 80 ns;
 
BEGIN
	UUT: ffms PORT MAP(
	Clk => Clk, 
	D => D, 
	Q => Q
   );
	
	  -- Clock process definitions
   Clk_process :process
   begin
		Clk <= '0';
		wait for Clk_period/2;
		Clk <= '1';
		wait for Clk_period/2;
   end process;
 



-- *** Test Bench - User Defined Section ***
   tb : PROCESS
   BEGIN
	
	D <= '0','1' after 180 ns,
	'0' after 220 ns, 
	'1' after 226 ns,
	'0' after 250 ns, '1' after 300 ns, '0' after 330 ns;
	
      WAIT; -- will wait forever
   END PROCESS;
-- *** End Test Bench - User Defined Section ***

END;
