----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    15:45:38 03/05/2019 
-- Design Name: 
-- Module Name:    XOR_Inversion - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity XOR_Inversion is
	generic( N: integer:= 8);
	Port ( 	
			input : in  STD_LOGIC_VECTOR (N - 1 downto 0);
         inverti : in  STD_LOGIC;
         output : out  STD_LOGIC_VECTOR (N - 1 downto 0));
end XOR_Inversion;

architecture Dataflow of XOR_Inversion is

signal temp :   STD_LOGIC_VECTOR (N - 1 downto 0);
begin
	XOR_Istanziation:for i in N-1 downto 0 generate
		temp(i)<=input(i) xor inverti;
	end generate XOR_Istanziation;
	output<= temp;


end Dataflow;

